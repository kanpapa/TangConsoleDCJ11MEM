parameter M=16;
parameter N=32;
parameter MSB=32;
parameter LATENCY=34;
